magic
tech sky130A
magscale 1 2
timestamp 1740548957
<< error_p >>
rect 6012 470 6132 490
rect 6656 470 6776 490
rect 8588 470 8708 490
rect 10520 470 10640 490
rect 11808 470 11928 490
rect 13648 470 13768 490
<< metal2 >>
rect 4066 40746 4122 41000
rect 3988 40718 4122 40746
rect 3988 40474 4016 40718
rect 4066 40600 4122 40718
rect 4710 40746 4766 41000
rect 5354 40746 5410 41000
rect 5998 40746 6054 41000
rect 6642 40746 6698 41000
rect 7286 40746 7342 41000
rect 7930 40746 7986 41000
rect 8574 40746 8630 41000
rect 9218 40746 9274 41000
rect 9862 40746 9918 41000
rect 10506 40746 10562 41000
rect 11150 40746 11206 41000
rect 11794 40746 11850 41000
rect 12438 40746 12494 41000
rect 13082 40746 13138 41000
rect 13726 40746 13782 41000
rect 14370 40746 14426 41000
rect 15014 40746 15070 41000
rect 4710 40718 4844 40746
rect 4710 40600 4766 40718
rect 3988 40446 4108 40474
rect 4080 40436 4108 40446
rect 4816 40436 4844 40718
rect 5354 40718 5488 40746
rect 5354 40600 5410 40718
rect 5460 40436 5488 40718
rect 5998 40718 6132 40746
rect 5998 40600 6054 40718
rect 6104 40436 6132 40718
rect 6642 40718 6776 40746
rect 6642 40600 6698 40718
rect 6748 40436 6776 40718
rect 7286 40718 7420 40746
rect 7286 40600 7342 40718
rect 7392 40436 7420 40718
rect 7930 40718 8064 40746
rect 7930 40600 7986 40718
rect 8036 40436 8064 40718
rect 8574 40718 8708 40746
rect 8574 40600 8630 40718
rect 8680 40436 8708 40718
rect 9218 40718 9352 40746
rect 9218 40600 9274 40718
rect 9324 40436 9352 40718
rect 9862 40718 9996 40746
rect 9862 40600 9918 40718
rect 9968 40436 9996 40718
rect 10506 40718 10640 40746
rect 10506 40600 10562 40718
rect 10612 40436 10640 40718
rect 11150 40718 11284 40746
rect 11150 40600 11206 40718
rect 11256 40436 11284 40718
rect 11794 40718 11928 40746
rect 11794 40600 11850 40718
rect 11900 40436 11928 40718
rect 12438 40718 12572 40746
rect 12438 40600 12494 40718
rect 12544 40436 12572 40718
rect 13082 40718 13216 40746
rect 13082 40600 13138 40718
rect 13188 40436 13216 40718
rect 13648 40718 13782 40746
rect 13648 40436 13676 40718
rect 13726 40600 13782 40718
rect 14108 40718 14426 40746
rect 14108 40436 14136 40718
rect 14370 40600 14426 40718
rect 14660 40718 15070 40746
rect 14660 40436 14688 40718
rect 15014 40600 15070 40718
rect 15566 40746 15622 40769
rect 15658 40746 15714 41000
rect 15566 40718 15714 40746
rect 15566 40695 15622 40718
rect 15658 40600 15714 40718
rect 16302 40746 16358 41000
rect 16946 40746 17002 41000
rect 17590 40746 17646 41000
rect 17682 40746 17738 40769
rect 16302 40718 16528 40746
rect 16302 40600 16358 40718
rect 16500 40436 16528 40718
rect 16946 40718 17080 40746
rect 16946 40600 17002 40718
rect 17052 40436 17080 40718
rect 17590 40718 17738 40746
rect 17590 40600 17646 40718
rect 17682 40695 17738 40718
rect 18234 40746 18290 41000
rect 18510 40746 18566 40769
rect 18234 40718 18566 40746
rect 18234 40600 18290 40718
rect 18510 40695 18566 40718
rect 18878 40746 18934 41000
rect 18878 40718 19012 40746
rect 18878 40600 18934 40718
rect 18984 40436 19012 40718
rect 19522 40600 19578 41000
rect 20166 40600 20222 41000
rect 20810 40600 20866 41000
rect 21454 40600 21510 41000
rect 22098 40600 22154 41000
rect 22742 40600 22798 41000
rect 23386 40600 23442 41000
rect 24030 40600 24086 41000
rect 24674 40746 24730 41000
rect 24412 40718 24730 40746
rect 24412 40436 24440 40718
rect 24674 40600 24730 40718
rect 25134 40746 25190 40769
rect 25318 40746 25374 41000
rect 25134 40718 25374 40746
rect 25134 40695 25190 40718
rect 25318 40600 25374 40718
rect 25870 40746 25926 40769
rect 25962 40746 26018 41000
rect 25870 40718 26018 40746
rect 25870 40695 25926 40718
rect 25962 40600 26018 40718
rect 26606 40600 26662 41000
rect 27250 40600 27306 41000
rect 27894 40600 27950 41000
rect 28538 40600 28594 41000
rect 29182 40600 29238 41000
rect 29826 40746 29882 41000
rect 30470 40746 30526 41000
rect 29826 40718 30144 40746
rect 29826 40600 29882 40718
rect 30116 40436 30144 40718
rect 30392 40718 30526 40746
rect 30392 40436 30420 40718
rect 30470 40600 30526 40718
rect 31114 40600 31170 41000
rect 2792 400 2820 470
rect 3436 400 3464 470
rect 4080 400 4108 470
rect 4724 400 4752 470
rect 5368 400 5396 470
rect 6012 462 6132 470
rect 6012 400 6040 462
rect 2778 0 2834 400
rect 3422 0 3478 400
rect 4066 0 4122 400
rect 4710 0 4766 400
rect 5354 0 5410 400
rect 5998 0 6054 400
rect 6104 202 6132 462
rect 6656 462 6776 470
rect 6656 400 6684 462
rect 6092 138 6144 202
rect 6642 0 6698 400
rect 6748 134 6776 462
rect 7300 400 7328 470
rect 7944 400 7972 470
rect 8588 462 8708 470
rect 8588 400 8616 462
rect 6736 70 6788 134
rect 7286 0 7342 400
rect 7930 0 7986 400
rect 8574 0 8630 400
rect 8680 66 8708 462
rect 9232 400 9260 470
rect 9876 400 9904 470
rect 10232 410 10284 470
rect 10520 462 10640 470
rect 10520 400 10548 462
rect 8668 2 8720 66
rect 9218 0 9274 400
rect 9862 0 9918 400
rect 10506 0 10562 400
rect 10612 105 10640 462
rect 11164 400 11192 470
rect 10598 31 10654 105
rect 11150 0 11206 400
rect 11348 202 11376 470
rect 11716 406 11744 470
rect 11808 462 11928 470
rect 11704 342 11756 406
rect 11808 400 11836 462
rect 11336 138 11388 202
rect 11794 0 11850 400
rect 11900 241 11928 462
rect 12452 400 12480 470
rect 13096 400 13124 470
rect 13188 406 13216 470
rect 13372 406 13400 470
rect 11886 167 11942 241
rect 12438 0 12494 400
rect 13082 0 13138 400
rect 13176 342 13228 406
rect 13360 342 13412 406
rect 13464 354 13492 470
rect 13648 462 13768 470
rect 13648 354 13676 462
rect 13740 400 13768 462
rect 14384 400 14412 470
rect 15028 400 15056 470
rect 15672 400 15700 470
rect 16316 400 16344 470
rect 16960 400 16988 470
rect 17604 400 17632 470
rect 13464 326 13676 354
rect 13726 0 13782 400
rect 14370 0 14426 400
rect 15014 0 15070 400
rect 15658 0 15714 400
rect 16302 0 16358 400
rect 16946 0 17002 400
rect 17590 0 17646 400
rect 18064 270 18092 470
rect 18248 400 18276 470
rect 18892 400 18920 470
rect 18052 206 18104 270
rect 18234 0 18290 400
rect 18878 0 18934 400
rect 18984 270 19012 470
rect 19536 400 19564 470
rect 20272 456 20300 470
rect 20180 428 20300 456
rect 20180 400 20208 428
rect 20824 400 20852 470
rect 18972 206 19024 270
rect 19522 0 19578 400
rect 20166 0 20222 400
rect 20810 0 20866 400
rect 21284 134 21312 470
rect 21468 400 21496 470
rect 21916 410 21968 470
rect 22112 400 22140 470
rect 22388 406 22416 470
rect 21272 70 21324 134
rect 21454 0 21510 400
rect 22098 0 22154 400
rect 22376 342 22428 406
rect 22756 400 22784 470
rect 22836 410 22888 470
rect 22742 0 22798 400
rect 22940 66 22968 470
rect 23400 400 23428 470
rect 22928 2 22980 66
rect 23386 0 23442 400
rect 23768 354 23796 470
rect 23952 428 24072 456
rect 23952 354 23980 428
rect 24044 400 24072 428
rect 23768 326 23980 354
rect 24030 0 24086 400
rect 24504 338 24532 470
rect 24688 400 24716 470
rect 25332 400 25360 470
rect 25976 400 26004 470
rect 26620 400 26648 470
rect 27264 400 27292 470
rect 27804 456 27856 470
rect 27804 428 27936 456
rect 27804 410 27856 428
rect 27908 400 27936 428
rect 24492 274 24544 338
rect 24674 0 24730 400
rect 25318 0 25374 400
rect 25962 0 26018 400
rect 26606 0 26662 400
rect 27250 0 27306 400
rect 27894 0 27950 400
rect 28000 241 28028 470
rect 28552 400 28580 470
rect 29196 400 29224 470
rect 29840 400 29868 470
rect 30484 400 30512 470
rect 27986 167 28042 241
rect 28538 0 28594 400
rect 29182 0 29238 400
rect 29826 0 29882 400
rect 30470 0 30526 400
rect 31036 270 31064 470
rect 31128 400 31156 470
rect 31024 206 31076 270
rect 31114 0 31170 400
<< labels >>
flabel metal2 s 11794 0 11850 400 0 FreeSans 280 90 0 0 B[0]
port 1 nsew
flabel metal2 s 5354 0 5410 400 0 FreeSans 280 90 0 0 B[10]
port 2 nsew
flabel metal2 s 4710 0 4766 400 0 FreeSans 280 90 0 0 B[11]
port 3 nsew
flabel metal2 s 11150 0 11206 400 0 FreeSans 280 90 0 0 B[1]
port 4 nsew
flabel metal2 s 10506 0 10562 400 0 FreeSans 280 90 0 0 B[2]
port 5 nsew
flabel metal2 s 9862 0 9918 400 0 FreeSans 280 90 0 0 B[3]
port 6 nsew
flabel metal2 s 9218 0 9274 400 0 FreeSans 280 90 0 0 B[4]
port 7 nsew
flabel metal2 s 8574 0 8630 400 0 FreeSans 280 90 0 0 B[5]
port 8 nsew
flabel metal2 s 7930 0 7986 400 0 FreeSans 280 90 0 0 B[6]
port 9 nsew
flabel metal2 s 7286 0 7342 400 0 FreeSans 280 90 0 0 B[7]
port 10 nsew
flabel metal2 s 6642 0 6698 400 0 FreeSans 280 90 0 0 B[8]
port 11 nsew
flabel metal2 s 5998 0 6054 400 0 FreeSans 280 90 0 0 B[9]
port 12 nsew
flabel metal2 s 4066 0 4122 400 0 FreeSans 280 90 0 0 Bvb[0]
port 13 nsew
flabel metal2 s 3422 0 3478 400 0 FreeSans 280 90 0 0 Bvb[1]
port 14 nsew
flabel metal2 s 2778 0 2834 400 0 FreeSans 280 90 0 0 Bvb[2]
port 15 nsew
flabel metal2 s 21454 0 21510 400 0 FreeSans 280 90 0 0 G[0]
port 16 nsew
flabel metal2 s 15014 0 15070 400 0 FreeSans 280 90 0 0 G[10]
port 17 nsew
flabel metal2 s 14370 0 14426 400 0 FreeSans 280 90 0 0 G[11]
port 18 nsew
flabel metal2 s 20810 0 20866 400 0 FreeSans 280 90 0 0 G[1]
port 19 nsew
flabel metal2 s 20166 0 20222 400 0 FreeSans 280 90 0 0 G[2]
port 20 nsew
flabel metal2 s 19522 0 19578 400 0 FreeSans 280 90 0 0 G[3]
port 21 nsew
flabel metal2 s 18878 0 18934 400 0 FreeSans 280 90 0 0 G[4]
port 22 nsew
flabel metal2 s 18234 0 18290 400 0 FreeSans 280 90 0 0 G[5]
port 23 nsew
flabel metal2 s 17590 0 17646 400 0 FreeSans 280 90 0 0 G[6]
port 24 nsew
flabel metal2 s 16946 0 17002 400 0 FreeSans 280 90 0 0 G[7]
port 25 nsew
flabel metal2 s 16302 0 16358 400 0 FreeSans 280 90 0 0 G[8]
port 26 nsew
flabel metal2 s 15658 0 15714 400 0 FreeSans 280 90 0 0 G[9]
port 27 nsew
flabel metal2 s 13726 0 13782 400 0 FreeSans 280 90 0 0 Gvb[0]
port 28 nsew
flabel metal2 s 13082 0 13138 400 0 FreeSans 280 90 0 0 Gvb[1]
port 29 nsew
flabel metal2 s 12438 0 12494 400 0 FreeSans 280 90 0 0 Gvb[2]
port 30 nsew
flabel metal2 s 31114 0 31170 400 0 FreeSans 280 90 0 0 R[0]
port 31 nsew
flabel metal2 s 24674 0 24730 400 0 FreeSans 280 90 0 0 R[10]
port 32 nsew
flabel metal2 s 24030 0 24086 400 0 FreeSans 280 90 0 0 R[11]
port 33 nsew
flabel metal2 s 30470 0 30526 400 0 FreeSans 280 90 0 0 R[1]
port 34 nsew
flabel metal2 s 29826 0 29882 400 0 FreeSans 280 90 0 0 R[2]
port 35 nsew
flabel metal2 s 29182 0 29238 400 0 FreeSans 280 90 0 0 R[3]
port 36 nsew
flabel metal2 s 28538 0 28594 400 0 FreeSans 280 90 0 0 R[4]
port 37 nsew
flabel metal2 s 27894 0 27950 400 0 FreeSans 280 90 0 0 R[5]
port 38 nsew
flabel metal2 s 27250 0 27306 400 0 FreeSans 280 90 0 0 R[6]
port 39 nsew
flabel metal2 s 26606 0 26662 400 0 FreeSans 280 90 0 0 R[7]
port 40 nsew
flabel metal2 s 25962 0 26018 400 0 FreeSans 280 90 0 0 R[8]
port 41 nsew
flabel metal2 s 25318 0 25374 400 0 FreeSans 280 90 0 0 R[9]
port 42 nsew
flabel metal2 s 23386 0 23442 400 0 FreeSans 280 90 0 0 Rvb[0]
port 43 nsew
flabel metal2 s 22742 0 22798 400 0 FreeSans 280 90 0 0 Rvb[1]
port 44 nsew
flabel metal2 s 22098 0 22154 400 0 FreeSans 280 90 0 0 Rvb[2]
port 45 nsew
flabel metal2 s 30470 40600 30526 41000 0 FreeSans 280 90 0 0 clk
port 48 nsew
flabel metal2 s 31114 40600 31170 41000 0 FreeSans 280 90 0 0 ena
port 49 nsew
flabel metal2 s 29826 40600 29882 41000 0 FreeSans 280 90 0 0 rst_n
port 50 nsew
flabel metal2 s 29182 40600 29238 41000 0 FreeSans 280 90 0 0 ui_in[0]
port 51 nsew
flabel metal2 s 28538 40600 28594 41000 0 FreeSans 280 90 0 0 ui_in[1]
port 52 nsew
flabel metal2 s 27894 40600 27950 41000 0 FreeSans 280 90 0 0 ui_in[2]
port 53 nsew
flabel metal2 s 27250 40600 27306 41000 0 FreeSans 280 90 0 0 ui_in[3]
port 54 nsew
flabel metal2 s 26606 40600 26662 41000 0 FreeSans 280 90 0 0 ui_in[4]
port 55 nsew
flabel metal2 s 25962 40600 26018 41000 0 FreeSans 280 90 0 0 ui_in[5]
port 56 nsew
flabel metal2 s 25318 40600 25374 41000 0 FreeSans 280 90 0 0 ui_in[6]
port 57 nsew
flabel metal2 s 24674 40600 24730 41000 0 FreeSans 280 90 0 0 ui_in[7]
port 58 nsew
flabel metal2 s 24030 40600 24086 41000 0 FreeSans 280 90 0 0 uio_in[0]
port 59 nsew
flabel metal2 s 23386 40600 23442 41000 0 FreeSans 280 90 0 0 uio_in[1]
port 60 nsew
flabel metal2 s 22742 40600 22798 41000 0 FreeSans 280 90 0 0 uio_in[2]
port 61 nsew
flabel metal2 s 22098 40600 22154 41000 0 FreeSans 280 90 0 0 uio_in[3]
port 62 nsew
flabel metal2 s 21454 40600 21510 41000 0 FreeSans 280 90 0 0 uio_in[4]
port 63 nsew
flabel metal2 s 20810 40600 20866 41000 0 FreeSans 280 90 0 0 uio_in[5]
port 64 nsew
flabel metal2 s 20166 40600 20222 41000 0 FreeSans 280 90 0 0 uio_in[6]
port 65 nsew
flabel metal2 s 19522 40600 19578 41000 0 FreeSans 280 90 0 0 uio_in[7]
port 66 nsew
flabel metal2 s 8574 40600 8630 41000 0 FreeSans 280 90 0 0 uio_oe[0]
port 67 nsew
flabel metal2 s 7930 40600 7986 41000 0 FreeSans 280 90 0 0 uio_oe[1]
port 68 nsew
flabel metal2 s 7286 40600 7342 41000 0 FreeSans 280 90 0 0 uio_oe[2]
port 69 nsew
flabel metal2 s 6642 40600 6698 41000 0 FreeSans 280 90 0 0 uio_oe[3]
port 70 nsew
flabel metal2 s 5998 40600 6054 41000 0 FreeSans 280 90 0 0 uio_oe[4]
port 71 nsew
flabel metal2 s 5354 40600 5410 41000 0 FreeSans 280 90 0 0 uio_oe[5]
port 72 nsew
flabel metal2 s 4710 40600 4766 41000 0 FreeSans 280 90 0 0 uio_oe[6]
port 73 nsew
flabel metal2 s 4066 40600 4122 41000 0 FreeSans 280 90 0 0 uio_oe[7]
port 74 nsew
flabel metal2 s 13726 40600 13782 41000 0 FreeSans 280 90 0 0 uio_out[0]
port 75 nsew
flabel metal2 s 13082 40600 13138 41000 0 FreeSans 280 90 0 0 uio_out[1]
port 76 nsew
flabel metal2 s 12438 40600 12494 41000 0 FreeSans 280 90 0 0 uio_out[2]
port 77 nsew
flabel metal2 s 11794 40600 11850 41000 0 FreeSans 280 90 0 0 uio_out[3]
port 78 nsew
flabel metal2 s 11150 40600 11206 41000 0 FreeSans 280 90 0 0 uio_out[4]
port 79 nsew
flabel metal2 s 10506 40600 10562 41000 0 FreeSans 280 90 0 0 uio_out[5]
port 80 nsew
flabel metal2 s 9862 40600 9918 41000 0 FreeSans 280 90 0 0 uio_out[6]
port 81 nsew
flabel metal2 s 9218 40600 9274 41000 0 FreeSans 280 90 0 0 uio_out[7]
port 82 nsew
flabel metal2 s 18878 40600 18934 41000 0 FreeSans 280 90 0 0 uo_out[0]
port 83 nsew
flabel metal2 s 18234 40600 18290 41000 0 FreeSans 280 90 0 0 uo_out[1]
port 84 nsew
flabel metal2 s 17590 40600 17646 41000 0 FreeSans 280 90 0 0 uo_out[2]
port 85 nsew
flabel metal2 s 16946 40600 17002 41000 0 FreeSans 280 90 0 0 uo_out[3]
port 86 nsew
flabel metal2 s 16302 40600 16358 41000 0 FreeSans 280 90 0 0 uo_out[4]
port 87 nsew
flabel metal2 s 15658 40600 15714 41000 0 FreeSans 280 90 0 0 uo_out[5]
port 88 nsew
flabel metal2 s 15014 40600 15070 41000 0 FreeSans 280 90 0 0 uo_out[6]
port 89 nsew
flabel metal2 s 14370 40600 14426 41000 0 FreeSans 280 90 0 0 uo_out[7]
port 90 nsew
<< properties >>
string FIXED_BBOX 0 0 63000 41000
<< end >>
